* D:\Archivos\Proyecto\Practica3.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 15 17:35:02 2019



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Practica3.net"
.INC "Practica3.als"


.probe


.END
