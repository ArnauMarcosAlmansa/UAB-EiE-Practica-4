* C:\Users\arnau\Desktop\repos\UAB-EiE-Practica-4\recursos\Ejercicio5.sch

* Schematics Version 9.1 - Web Update 1
* Mon Oct 21 13:49:50 2019



** Analysis setup **
.tran 0ns 0.04s
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ejercicio5.net"
.INC "Ejercicio5.als"


.probe


.END
