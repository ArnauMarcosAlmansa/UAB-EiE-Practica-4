* D:\Archivos\Proyecto\Ejercicio5.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 15 19:01:50 2019



** Analysis setup **
.tran 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ejercicio5.net"
.INC "Ejercicio5.als"


.probe


.END
